magic
tech sky130A
magscale 1 2
timestamp 1729215025
<< nwell >>
rect -177 -2062 822 995
<< nsubdiff >>
rect -141 925 -81 959
rect 726 925 786 959
rect -141 899 -107 925
rect 752 899 786 925
rect -141 -1992 -107 -1966
rect 752 -1992 786 -1966
rect -141 -2026 -81 -1992
rect 726 -2026 786 -1992
<< nsubdiffcont >>
rect -81 925 726 959
rect -141 -1966 -107 899
rect 752 -1966 786 899
rect -81 -2026 726 -1992
<< poly >>
rect -56 887 36 903
rect -56 853 -40 887
rect -6 853 36 887
rect -56 837 36 853
rect 6 804 36 837
rect 610 887 702 903
rect 610 853 652 887
rect 686 853 702 887
rect 610 837 702 853
rect 610 829 640 837
rect -57 107 35 123
rect 92 116 294 308
rect -57 73 -41 107
rect -7 73 35 107
rect -57 57 35 73
rect 5 24 35 57
rect 609 107 701 123
rect 609 73 651 107
rect 685 73 701 107
rect 609 57 701 73
rect 609 24 639 57
rect 94 -624 552 -470
rect 5 -1149 35 -1116
rect -57 -1165 35 -1149
rect -57 -1199 -41 -1165
rect -7 -1199 35 -1165
rect -57 -1215 35 -1199
rect 609 -1151 639 -1118
rect 609 -1167 701 -1151
rect 609 -1201 651 -1167
rect 685 -1201 701 -1167
rect 352 -1378 550 -1212
rect 609 -1217 701 -1201
rect 5 -1904 35 -1871
rect -57 -1920 35 -1904
rect -57 -1954 -41 -1920
rect -7 -1954 35 -1920
rect -57 -1970 35 -1954
rect 609 -1904 639 -1873
rect 609 -1920 701 -1904
rect 609 -1954 651 -1920
rect 685 -1954 701 -1920
rect 609 -1970 701 -1954
<< polycont >>
rect -40 853 -6 887
rect 652 853 686 887
rect -41 73 -7 107
rect 651 73 685 107
rect -41 -1199 -7 -1165
rect 651 -1201 685 -1167
rect -41 -1954 -7 -1920
rect 651 -1954 685 -1920
<< locali >>
rect -141 925 -81 959
rect 726 925 786 959
rect -141 899 -107 925
rect 752 899 786 925
rect -56 853 -40 887
rect -6 853 10 887
rect 636 853 652 887
rect 686 853 702 887
rect -40 804 -6 853
rect 652 802 686 853
rect -57 73 -41 107
rect -7 73 9 107
rect 635 73 651 107
rect 685 73 701 107
rect -41 24 -7 73
rect 651 24 685 73
rect -41 -1165 -7 -1116
rect -57 -1199 -41 -1165
rect -7 -1199 9 -1165
rect 651 -1167 685 -1118
rect 635 -1201 651 -1167
rect 685 -1201 701 -1167
rect -41 -1920 -7 -1871
rect 651 -1920 685 -1873
rect -57 -1954 -41 -1920
rect -7 -1954 9 -1920
rect 635 -1954 651 -1920
rect 685 -1954 701 -1920
rect -141 -1992 -107 -1966
rect 752 -1992 786 -1966
rect -141 -2026 -81 -1992
rect 726 -2026 786 -1992
<< viali >>
rect 653 925 687 959
rect -40 853 -6 887
rect 652 853 686 887
rect -41 73 -7 107
rect 651 73 685 107
rect -41 -1199 -7 -1165
rect 651 -1201 685 -1167
rect -41 -1954 -7 -1920
rect 651 -1954 685 -1920
rect -41 -2026 -7 -1992
<< metal1 >>
rect 641 959 699 965
rect 641 931 653 959
rect 640 925 653 931
rect 687 925 699 959
rect 640 919 699 925
rect -52 887 6 893
rect -52 853 -40 887
rect -6 853 6 887
rect -52 847 6 853
rect 640 887 698 919
rect 640 853 652 887
rect 686 853 698 887
rect 640 847 698 853
rect -46 804 0 847
rect 646 805 692 847
rect -48 793 87 803
rect -58 416 -48 793
rect 4 416 87 793
rect -48 403 87 416
rect 299 363 346 804
rect 558 405 693 805
rect 558 363 604 405
rect 299 317 386 363
rect 513 317 604 363
rect -53 107 5 113
rect -53 73 -41 107
rect -7 73 5 107
rect -53 67 5 73
rect -47 24 -1 67
rect -46 -374 39 24
rect 92 -374 102 24
rect -46 -376 89 -374
rect 81 -632 123 -631
rect 32 -678 125 -632
rect 32 -723 101 -678
rect -51 -730 101 -723
rect -51 -1107 38 -730
rect 90 -749 101 -730
rect 90 -1107 100 -749
rect -51 -1109 99 -1107
rect -47 -1159 -1 -1116
rect 32 -1119 96 -1109
rect -53 -1165 5 -1159
rect -53 -1199 -41 -1165
rect -7 -1199 5 -1165
rect -53 -1205 5 -1199
rect 299 -1386 346 317
rect 639 107 697 113
rect 639 73 651 107
rect 685 73 697 107
rect 639 67 697 73
rect 548 23 612 25
rect 645 24 691 67
rect 548 13 691 23
rect 544 -364 554 13
rect 606 -364 691 13
rect 548 -377 691 -364
rect 548 -410 616 -377
rect 548 -417 613 -410
rect 515 -463 613 -417
rect 557 -724 692 -717
rect 539 -1118 549 -724
rect 606 -1117 692 -724
rect 606 -1118 616 -1117
rect 645 -1161 691 -1118
rect 639 -1167 697 -1161
rect 639 -1201 651 -1167
rect 685 -1201 697 -1167
rect 639 -1207 697 -1201
rect 41 -1432 130 -1386
rect 262 -1432 346 -1386
rect 41 -1473 87 -1432
rect -47 -1873 88 -1473
rect 299 -1872 346 -1432
rect 465 -1433 522 -1386
rect 557 -1485 692 -1472
rect 557 -1861 642 -1485
rect 694 -1861 704 -1485
rect 557 -1872 692 -1861
rect -47 -1914 -1 -1873
rect 645 -1914 691 -1873
rect -53 -1920 5 -1914
rect -53 -1954 -41 -1920
rect -7 -1954 5 -1920
rect -53 -1992 5 -1954
rect 639 -1920 697 -1914
rect 639 -1954 651 -1920
rect 685 -1954 697 -1920
rect 639 -1960 697 -1954
rect -53 -2026 -41 -1992
rect -7 -2026 5 -1992
rect -53 -2032 5 -2026
<< via1 >>
rect -48 416 4 793
rect 39 -374 92 24
rect 38 -1107 90 -730
rect 554 -364 606 13
rect 549 -1118 606 -724
rect 642 -1861 694 -1485
<< metal2 >>
rect -48 793 4 803
rect -49 416 -48 619
rect -49 406 4 416
rect -49 249 3 406
rect -56 239 4 249
rect -56 164 4 174
rect 640 235 696 245
rect 640 169 696 179
rect -53 -1235 2 164
rect 39 24 92 34
rect 554 22 606 23
rect 39 -384 92 -374
rect 552 13 608 22
rect 552 -39 554 13
rect 606 -39 608 13
rect 552 -375 608 -365
rect 40 -494 84 -384
rect 40 -600 601 -494
rect 40 -601 84 -600
rect 558 -714 600 -600
rect 36 -730 92 -720
rect 36 -1117 92 -1107
rect 549 -724 606 -714
rect 549 -1128 606 -1118
rect 642 -1231 694 169
rect -54 -1245 2 -1235
rect -54 -1311 2 -1301
rect 640 -1241 696 -1231
rect 640 -1313 696 -1303
rect 642 -1485 694 -1313
rect 642 -1871 694 -1861
<< via2 >>
rect -56 174 4 239
rect 640 179 696 235
rect 552 -364 554 -39
rect 554 -364 606 -39
rect 606 -364 608 -39
rect 552 -365 608 -364
rect 36 -1107 38 -730
rect 38 -1107 90 -730
rect 90 -1107 92 -730
rect -54 -1301 2 -1245
rect 640 -1303 696 -1241
<< metal3 >>
rect -66 240 14 244
rect -66 239 706 240
rect -66 174 -56 239
rect 4 235 706 239
rect 4 179 640 235
rect 696 179 706 235
rect 4 174 706 179
rect -66 169 14 174
rect 544 -39 618 -14
rect 544 -365 552 -39
rect 608 -365 618 -39
rect 544 -368 618 -365
rect 544 -513 619 -368
rect 25 -574 619 -513
rect 25 -727 102 -574
rect 26 -730 102 -727
rect 26 -1107 36 -730
rect 92 -1107 102 -730
rect 26 -1112 102 -1107
rect -64 -1241 12 -1240
rect 630 -1241 706 -1236
rect -64 -1245 640 -1241
rect -64 -1301 -54 -1245
rect 2 -1301 640 -1245
rect -64 -1302 640 -1301
rect -64 -1306 12 -1302
rect 630 -1303 640 -1302
rect 696 -1303 706 -1241
rect 630 -1308 706 -1303
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729133377
transform 1 0 20 0 1 -176
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729133377
transform 1 0 21 0 1 604
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729133377
transform 1 0 625 0 1 604
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729133377
transform 1 0 624 0 1 -176
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729133377
transform 1 0 624 0 1 -918
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729133377
transform 1 0 624 0 1 -1673
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729133377
transform 1 0 20 0 1 -918
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729133377
transform 1 0 20 0 1 -1673
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729147051
transform 1 0 323 0 1 604
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729147051
transform 1 0 322 0 1 -176
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729147051
transform 1 0 322 0 1 -918
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729147051
transform 1 0 322 0 1 -1673
box -323 -300 323 300
<< labels >>
flabel metal1 666 912 666 912 0 FreeSans 800 0 0 0 vdd
port 0 nsew
flabel metal2 666 -610 666 -610 0 FreeSans 800 0 0 0 d5
port 3 nsew
flabel metal3 573 -480 573 -480 0 FreeSans 800 0 0 0 d1
port 2 nsew
flabel metal2 59 -452 59 -452 0 FreeSans 800 0 0 0 d2
port 4 nsew
<< end >>
