magic
tech sky130A
magscale 1 2
timestamp 1729359112
<< viali >>
rect -307 2835 -249 2888
<< metal1 >>
rect -319 2888 -237 2894
rect -319 2835 -307 2888
rect -249 2835 819 2888
rect -319 2829 -237 2835
rect -307 1795 -249 2829
rect 761 2704 819 2835
rect 58 2107 68 2163
rect 124 2107 134 2163
rect 1469 2110 1479 2162
rect 1531 2110 1541 2162
rect -79 1369 -69 1421
rect -17 1409 -7 1421
rect 589 1409 617 1789
rect 1480 1596 1490 1648
rect 1542 1596 1552 1648
rect -17 1381 617 1409
rect 879 1397 889 1449
rect 941 1397 951 1449
rect -17 1369 -7 1381
rect -76 1105 -66 1157
rect -14 1154 -4 1157
rect -14 1109 288 1154
rect -14 1105 -4 1109
rect 892 -109 938 -16
rect 1040 -109 1050 -103
rect 892 -150 1050 -109
rect 892 -229 938 -150
rect 1040 -155 1050 -150
rect 1102 -155 1112 -103
rect 1557 -116 1567 -111
rect 1216 -159 1567 -116
rect 892 -263 999 -229
rect 1216 -417 1262 -159
rect 1557 -163 1567 -159
rect 1619 -163 1629 -111
<< via1 >>
rect 68 2107 124 2163
rect 1479 2110 1531 2162
rect -69 1369 -17 1421
rect 1490 1596 1542 1648
rect 889 1397 941 1449
rect -66 1105 -14 1157
rect 1050 -155 1102 -103
rect 1567 -163 1619 -111
<< metal2 >>
rect 972 2587 1024 2597
rect 68 2163 124 2173
rect 1479 2169 1531 2172
rect 68 2097 124 2107
rect 967 2162 1538 2169
rect 967 2110 1479 2162
rect 1531 2110 1538 2162
rect 967 2104 1538 2110
rect 1479 2100 1531 2104
rect 1490 1648 1542 1658
rect 1046 1596 1490 1648
rect 1490 1586 1542 1596
rect 889 1449 941 1459
rect -71 1423 -15 1433
rect -71 1357 -15 1367
rect 889 1199 941 1397
rect -66 1157 -14 1167
rect -909 1109 -66 1155
rect -909 848 -855 1109
rect -66 1095 -14 1105
rect 1050 -103 1102 -93
rect 1050 -165 1102 -155
rect 1496 -696 1532 1586
rect 1565 -109 1621 -99
rect 1565 -175 1621 -165
rect 1214 -744 1532 -696
<< via2 >>
rect 68 2107 124 2163
rect -71 1421 -15 1423
rect -71 1369 -69 1421
rect -69 1369 -17 1421
rect -17 1369 -15 1421
rect -71 1367 -15 1369
rect 1565 -111 1621 -109
rect 1565 -163 1567 -111
rect 1567 -163 1619 -111
rect 1619 -163 1621 -111
rect 1565 -165 1621 -163
<< metal3 >>
rect 56 2163 490 2174
rect 56 2107 68 2163
rect 124 2107 490 2163
rect 56 2096 490 2107
rect 1230 1729 1631 1791
rect -81 1423 -5 1428
rect -81 1367 -71 1423
rect -15 1367 -5 1423
rect -81 1075 -5 1367
rect -248 1009 -5 1075
rect 7 648 465 708
rect 7 322 67 648
rect -398 262 67 322
rect 1555 -109 1631 1729
rect 1555 -165 1565 -109
rect 1621 -165 1631 -109
rect 1555 -170 1631 -165
use NMOS  NMOS_0
timestamp 1729225705
transform 1 0 457 0 1 720
box -303 -743 1033 647
use NMOS_2  NMOS_2_0
timestamp 1729338435
transform 1 0 338 0 1 -670
box -184 -549 1124 447
use PMOS  PMOS_0
timestamp 1729215025
transform 1 0 -948 0 1 835
box -177 -2062 822 995
use PMOS_2  PMOS_2_0
timestamp 1729351298
transform 1 0 542 0 1 4469
box -388 -2963 853 -1702
<< labels >>
flabel viali -278 2859 -278 2859 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel via1 1505 2135 1505 2135 0 FreeSans 320 0 0 0 VIN
port 1 nsew
flabel via2 96 2135 96 2135 0 FreeSans 320 0 0 0 VIP
port 2 nsew
flabel via1 915 1423 915 1423 0 FreeSans 320 0 0 0 RS
port 3 nsew
flabel via1 1077 -129 1077 -129 0 FreeSans 320 0 0 0 GND
port 4 nsew
flabel via1 1516 1623 1516 1623 0 FreeSans 320 0 0 0 OUT
port 5 nsew
<< end >>
