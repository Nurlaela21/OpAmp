magic
tech sky130A
magscale 1 2
timestamp 1729351298
<< nwell >>
rect -388 -2963 853 -1702
<< nsubdiff >>
rect -352 -1772 -292 -1738
rect 757 -1772 817 -1738
rect -352 -1798 -318 -1772
rect 783 -1798 817 -1772
rect -352 -2893 -318 -2867
rect 783 -2893 817 -2867
rect -352 -2927 -292 -2893
rect 757 -2927 817 -2893
<< nsubdiffcont >>
rect -292 -1772 757 -1738
rect -352 -2867 -318 -1798
rect 783 -2867 817 -1798
rect -292 -2927 757 -2893
<< poly >>
rect -156 -2224 -126 -2198
rect -218 -2240 -126 -2224
rect -218 -2274 -202 -2240
rect -168 -2274 -126 -2240
rect -218 -2290 -126 -2274
rect 564 -2224 594 -2198
rect 564 -2240 656 -2224
rect 564 -2274 606 -2240
rect 640 -2274 656 -2240
rect 564 -2290 656 -2274
rect -218 -2391 -126 -2375
rect -218 -2425 -202 -2391
rect -168 -2425 -126 -2391
rect -218 -2441 -126 -2425
rect -156 -2467 -126 -2441
rect 564 -2391 656 -2375
rect 564 -2425 606 -2391
rect 640 -2425 656 -2391
rect 564 -2441 656 -2425
rect 564 -2467 594 -2441
<< polycont >>
rect -202 -2274 -168 -2240
rect 606 -2274 640 -2240
rect -202 -2425 -168 -2391
rect 606 -2425 640 -2391
<< locali >>
rect -352 -1772 -292 -1738
rect 757 -1772 817 -1738
rect -352 -1798 -318 -1772
rect 783 -1798 817 -1772
rect -218 -2274 -202 -2240
rect -168 -2274 -152 -2240
rect 590 -2274 606 -2240
rect 640 -2274 656 -2240
rect -218 -2425 -202 -2391
rect -168 -2425 -152 -2391
rect 590 -2425 606 -2391
rect 640 -2425 656 -2391
rect -352 -2893 -318 -2867
rect 783 -2893 817 -2867
rect -352 -2927 -292 -2893
rect 757 -2927 817 -2893
<< viali >>
rect 90 -1772 348 -1738
rect -202 -2274 -168 -2240
rect 606 -2274 640 -2240
rect -202 -2425 -168 -2391
rect 606 -2425 640 -2391
<< metal1 >>
rect 78 -1738 360 -1732
rect 78 -1772 90 -1738
rect 348 -1772 360 -1738
rect 78 -1778 360 -1772
rect -54 -1934 -44 -1882
rect 8 -1934 18 -1882
rect 104 -1934 113 -1882
rect 165 -1934 176 -1882
rect 262 -1934 273 -1882
rect 325 -1934 334 -1882
rect 420 -1934 430 -1882
rect 482 -1934 492 -1882
rect 193 -1984 245 -1974
rect -202 -2160 -123 -1984
rect -71 -2160 -61 -1984
rect -202 -2234 -168 -2160
rect -214 -2240 -156 -2234
rect -214 -2274 -202 -2240
rect -168 -2274 -156 -2240
rect -54 -2262 -44 -2210
rect 8 -2262 18 -2210
rect -214 -2280 -156 -2274
rect 46 -2308 76 -2151
rect 183 -2160 193 -1984
rect 245 -2160 255 -1984
rect 104 -2262 114 -2210
rect 166 -2262 176 -2210
rect 262 -2262 272 -2210
rect 324 -2262 334 -2210
rect 362 -2308 392 -2149
rect 499 -2160 509 -1984
rect 561 -2160 640 -1984
rect 420 -2262 430 -2210
rect 482 -2262 492 -2210
rect 606 -2234 640 -2160
rect 594 -2240 652 -2234
rect 594 -2274 606 -2240
rect 640 -2274 652 -2240
rect 594 -2280 652 -2274
rect 46 -2357 392 -2308
rect -214 -2391 -156 -2385
rect -214 -2425 -202 -2391
rect -168 -2425 -156 -2391
rect -214 -2431 -156 -2425
rect -202 -2500 -168 -2431
rect -54 -2455 -44 -2403
rect 8 -2455 18 -2403
rect -202 -2681 -123 -2505
rect -71 -2681 -61 -2505
rect 46 -2514 76 -2357
rect 104 -2455 114 -2403
rect 166 -2455 176 -2403
rect 262 -2455 272 -2403
rect 324 -2455 334 -2403
rect 183 -2681 193 -2505
rect 245 -2681 255 -2505
rect 362 -2512 392 -2357
rect 594 -2391 652 -2385
rect 420 -2455 430 -2403
rect 482 -2455 492 -2403
rect 594 -2425 606 -2391
rect 640 -2425 652 -2391
rect 594 -2431 652 -2425
rect 606 -2505 640 -2431
rect 499 -2681 509 -2505
rect 561 -2681 640 -2505
rect -55 -2783 -43 -2731
rect 9 -2783 17 -2731
rect 104 -2783 114 -2731
rect 166 -2783 176 -2731
rect 262 -2783 272 -2731
rect 324 -2783 334 -2731
rect 414 -2783 424 -2727
rect 480 -2783 490 -2727
<< via1 >>
rect -44 -1934 8 -1882
rect 113 -1934 165 -1882
rect 273 -1934 325 -1882
rect 430 -1934 482 -1882
rect -123 -2160 -71 -1984
rect -44 -2262 8 -2210
rect 193 -2160 245 -1984
rect 114 -2262 166 -2210
rect 272 -2262 324 -2210
rect 509 -2160 561 -1984
rect 430 -2262 482 -2210
rect -44 -2455 8 -2403
rect -123 -2681 -71 -2505
rect 114 -2455 166 -2403
rect 272 -2455 324 -2403
rect 193 -2681 245 -2505
rect 430 -2455 482 -2403
rect 509 -2681 561 -2505
rect -43 -2783 9 -2731
rect 114 -2783 166 -2731
rect 272 -2783 324 -2731
rect 424 -2783 480 -2727
<< metal2 >>
rect -288 -1844 245 -1792
rect -288 -2821 -244 -1844
rect -44 -1882 8 -1872
rect -44 -1944 8 -1934
rect 113 -1882 165 -1872
rect 113 -1944 165 -1934
rect -125 -1984 -69 -1974
rect -125 -2170 -69 -2160
rect 193 -1984 245 -1844
rect 273 -1882 325 -1872
rect 273 -1944 325 -1934
rect 430 -1882 482 -1872
rect 430 -1944 482 -1934
rect 193 -2170 245 -2160
rect 507 -1984 563 -1974
rect 507 -2170 563 -2160
rect -44 -2210 8 -2200
rect -44 -2300 8 -2262
rect 112 -2205 168 -2195
rect 112 -2262 114 -2261
rect 166 -2262 168 -2261
rect 112 -2271 168 -2262
rect 270 -2206 326 -2196
rect 114 -2272 166 -2271
rect 270 -2272 326 -2262
rect 430 -2210 482 -2200
rect 430 -2300 482 -2262
rect -44 -2365 482 -2300
rect -44 -2397 8 -2393
rect -46 -2403 10 -2397
rect -46 -2407 -44 -2403
rect 8 -2407 10 -2403
rect -46 -2473 10 -2463
rect 114 -2403 166 -2365
rect 114 -2465 166 -2455
rect 272 -2403 324 -2365
rect 272 -2465 324 -2455
rect 428 -2403 484 -2393
rect 428 -2469 484 -2459
rect -123 -2505 -71 -2495
rect -123 -2821 -71 -2681
rect 191 -2505 247 -2495
rect 191 -2691 247 -2681
rect 509 -2505 561 -2495
rect -43 -2731 9 -2721
rect -43 -2793 9 -2783
rect 114 -2731 166 -2721
rect 114 -2793 166 -2783
rect 272 -2731 324 -2721
rect 272 -2793 324 -2783
rect 424 -2727 480 -2717
rect 424 -2793 480 -2783
rect 509 -2821 561 -2681
rect -288 -2873 561 -2821
<< via2 >>
rect -125 -2160 -123 -1984
rect -123 -2160 -71 -1984
rect -71 -2160 -69 -1984
rect 507 -2160 509 -1984
rect 509 -2160 561 -1984
rect 561 -2160 563 -1984
rect 112 -2210 168 -2205
rect 112 -2261 114 -2210
rect 114 -2261 166 -2210
rect 166 -2261 168 -2210
rect 270 -2210 326 -2206
rect 270 -2262 272 -2210
rect 272 -2262 324 -2210
rect 324 -2262 326 -2210
rect -46 -2455 -44 -2407
rect -44 -2455 8 -2407
rect 8 -2455 10 -2407
rect -46 -2463 10 -2455
rect 428 -2455 430 -2403
rect 430 -2455 482 -2403
rect 482 -2455 484 -2403
rect 428 -2459 484 -2455
rect 191 -2681 193 -2505
rect 193 -2681 245 -2505
rect 245 -2681 247 -2505
<< metal3 >>
rect -135 -1869 751 -1808
rect -135 -1984 -59 -1869
rect -135 -2160 -125 -1984
rect -69 -2160 -59 -1984
rect -135 -2165 -59 -2160
rect 497 -1984 573 -1869
rect 497 -2160 507 -1984
rect 563 -2160 573 -1984
rect 497 -2165 573 -2160
rect 102 -2205 178 -2200
rect 102 -2261 112 -2205
rect 168 -2261 178 -2205
rect 102 -2295 178 -2261
rect 260 -2206 336 -2201
rect 260 -2262 270 -2206
rect 326 -2262 336 -2206
rect 260 -2295 336 -2262
rect -56 -2373 494 -2295
rect -56 -2407 20 -2373
rect -56 -2463 -46 -2407
rect 10 -2463 20 -2407
rect -56 -2468 20 -2463
rect 418 -2403 494 -2373
rect 418 -2459 428 -2403
rect 484 -2459 494 -2403
rect 418 -2464 494 -2459
rect 181 -2505 257 -2500
rect 181 -2681 191 -2505
rect 247 -2681 257 -2505
rect 181 -2797 257 -2681
rect 688 -2797 751 -1869
rect 181 -2858 751 -2797
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729348687
transform 1 0 579 0 1 -2072
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729348687
transform 1 0 -141 0 1 -2072
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729348687
transform 1 0 -141 0 1 -2593
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729348687
transform 1 0 579 0 1 -2593
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_V8EW5L  sky130_fd_pr__pfet_01v8_V8EW5L_0
timestamp 1729344401
transform 1 0 219 0 1 -2593
box -381 -200 381 200
use sky130_fd_pr__pfet_01v8_V8EW5L  sky130_fd_pr__pfet_01v8_V8EW5L_1
timestamp 1729344401
transform 1 0 219 0 1 -2072
box -381 -200 381 200
<< labels >>
flabel viali 227 -1755 227 -1755 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal1 376 -2240 376 -2240 0 FreeSans 800 0 0 0 D5
port 1 nsew
flabel metal3 712 -1846 712 -1846 0 FreeSans 800 0 0 0 D6
port 4 nsew
flabel metal2 -260 -2848 -260 -2848 0 FreeSans 800 0 0 0 OUT
port 5 nsew
flabel metal2 302 -2383 302 -2383 0 FreeSans 800 0 0 0 VIN
port 7 nsew
flabel metal3 140 -2277 140 -2277 0 FreeSans 800 0 0 0 VIP
port 8 nsew
<< end >>
